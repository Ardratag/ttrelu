VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_ardratag_tt_relu
  CLASS BLOCK ;
  FOREIGN tt_um_ardratag_tt_relu ;
  ORIGIN -1.000 0.000 ;
  SIZE 157.850 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 66.450 9.840 68.520 11.460 ;
        RECT 133.330 9.520 135.400 11.140 ;
      LAYER li1 ;
        RECT 90.150 13.925 90.990 13.930 ;
        RECT 67.230 13.345 90.990 13.925 ;
        RECT 67.230 11.760 67.590 13.345 ;
        RECT 67.820 11.760 68.160 11.860 ;
        RECT 67.230 11.580 68.160 11.760 ;
        RECT 67.230 11.150 67.400 11.580 ;
        RECT 67.820 11.510 68.160 11.580 ;
        RECT 66.630 10.150 67.400 11.150 ;
        RECT 67.230 8.470 67.400 10.150 ;
        RECT 67.670 10.130 67.840 11.170 ;
        RECT 67.670 8.470 67.840 9.510 ;
        RECT 68.110 9.490 68.280 11.170 ;
        RECT 68.110 8.490 68.780 9.490 ;
        RECT 64.380 7.960 67.710 8.060 ;
        RECT 68.110 7.960 68.280 8.490 ;
        RECT 64.380 7.790 68.280 7.960 ;
        RECT 64.380 7.700 67.710 7.790 ;
        RECT 64.380 2.040 64.840 7.700 ;
        RECT 90.150 2.590 90.990 13.345 ;
        RECT 134.110 11.750 157.130 12.280 ;
        RECT 134.110 11.440 134.530 11.750 ;
        RECT 134.700 11.440 135.040 11.540 ;
        RECT 134.110 11.270 135.040 11.440 ;
        RECT 134.110 10.830 134.280 11.270 ;
        RECT 134.700 11.190 135.040 11.270 ;
        RECT 133.510 9.830 134.280 10.830 ;
        RECT 134.110 8.150 134.280 9.830 ;
        RECT 134.550 9.810 134.720 10.850 ;
        RECT 134.550 8.150 134.720 9.190 ;
        RECT 134.990 9.170 135.160 10.850 ;
        RECT 134.990 8.170 135.660 9.170 ;
        RECT 112.120 7.640 130.480 7.660 ;
        RECT 134.240 7.640 134.590 7.740 ;
        RECT 134.990 7.640 135.160 8.170 ;
        RECT 112.120 7.480 135.160 7.640 ;
        RECT 112.120 7.470 122.990 7.480 ;
        RECT 128.160 7.470 135.160 7.480 ;
        RECT 112.120 7.430 113.200 7.470 ;
        RECT 112.120 2.850 113.190 7.430 ;
        RECT 134.240 7.380 134.590 7.470 ;
        RECT 156.550 5.460 157.130 11.750 ;
        RECT 156.140 4.650 157.460 5.460 ;
        RECT 45.750 1.070 64.840 2.040 ;
        RECT 89.590 1.280 91.650 2.590 ;
        RECT 111.600 1.470 113.850 2.850 ;
      LAYER mcon ;
        RECT 67.230 10.210 67.400 11.090 ;
        RECT 67.670 10.210 67.840 11.090 ;
        RECT 68.110 10.210 68.280 11.090 ;
        RECT 67.230 8.550 67.400 9.430 ;
        RECT 67.670 8.550 67.840 9.430 ;
        RECT 68.110 8.550 68.280 9.430 ;
        RECT 134.110 9.890 134.280 10.770 ;
        RECT 134.550 9.890 134.720 10.770 ;
        RECT 134.990 9.890 135.160 10.770 ;
        RECT 134.110 8.230 134.280 9.110 ;
        RECT 134.550 8.230 134.720 9.110 ;
        RECT 134.990 8.230 135.160 9.110 ;
        RECT 156.530 4.830 157.110 5.320 ;
        RECT 46.090 1.270 46.800 1.900 ;
        RECT 89.890 1.570 91.220 2.360 ;
        RECT 112.120 1.720 113.170 2.570 ;
      LAYER met1 ;
        RECT 67.200 10.150 67.430 11.150 ;
        RECT 67.640 9.800 67.870 11.150 ;
        RECT 68.080 10.150 68.310 11.150 ;
        RECT 134.080 9.830 134.310 10.830 ;
        RECT 67.640 9.660 69.930 9.800 ;
        RECT 67.200 8.490 67.430 9.490 ;
        RECT 67.640 8.490 67.870 9.490 ;
        RECT 68.080 8.490 68.310 9.490 ;
        RECT 69.650 6.650 69.930 9.660 ;
        RECT 134.520 9.480 134.750 10.830 ;
        RECT 134.960 9.830 135.190 10.830 ;
        RECT 134.520 9.340 136.300 9.480 ;
        RECT 134.080 8.170 134.310 9.170 ;
        RECT 134.520 8.170 134.750 9.170 ;
        RECT 134.960 8.170 135.190 9.170 ;
        RECT 136.030 6.690 136.300 9.340 ;
        RECT 68.150 6.320 69.930 6.650 ;
        RECT 134.470 6.350 136.300 6.690 ;
        RECT 68.150 2.570 68.880 6.320 ;
        RECT 68.150 2.560 68.950 2.570 ;
        RECT 45.750 1.070 47.180 2.040 ;
        RECT 67.740 1.500 69.320 2.560 ;
        RECT 89.590 1.280 91.650 2.590 ;
        RECT 111.600 1.470 113.850 2.850 ;
        RECT 134.470 2.800 135.060 6.350 ;
        RECT 156.140 4.650 157.460 5.460 ;
        RECT 134.110 1.700 135.430 2.800 ;
      LAYER via ;
        RECT 46.090 1.270 46.800 1.900 ;
        RECT 68.150 1.690 68.890 2.410 ;
        RECT 89.890 1.570 91.220 2.360 ;
        RECT 156.530 4.830 157.110 5.320 ;
        RECT 112.120 1.720 113.170 2.570 ;
        RECT 134.470 2.010 135.070 2.570 ;
      LAYER met2 ;
        RECT 156.140 4.650 157.460 5.460 ;
        RECT 45.750 1.070 47.180 2.040 ;
        RECT 67.740 1.500 69.320 2.560 ;
        RECT 89.590 1.280 91.650 2.590 ;
        RECT 111.600 1.470 113.850 2.850 ;
        RECT 134.110 1.700 135.430 2.800 ;
      LAYER via2 ;
        RECT 156.530 4.830 157.110 5.320 ;
        RECT 46.090 1.270 46.800 1.900 ;
        RECT 68.150 1.690 68.890 2.410 ;
        RECT 89.890 1.570 91.220 2.360 ;
        RECT 112.120 1.720 113.170 2.570 ;
        RECT 134.470 2.010 135.070 2.570 ;
      LAYER met3 ;
        RECT 156.140 4.650 157.460 5.460 ;
        RECT 45.750 1.070 47.180 2.040 ;
        RECT 67.740 1.500 69.320 2.560 ;
        RECT 89.590 1.280 91.650 2.590 ;
        RECT 111.600 1.470 113.850 2.850 ;
        RECT 134.110 1.700 135.430 2.800 ;
      LAYER via3 ;
        RECT 156.530 4.830 157.110 5.320 ;
        RECT 46.090 1.270 46.800 1.900 ;
        RECT 68.150 1.690 68.890 2.410 ;
        RECT 89.890 1.570 91.220 2.360 ;
        RECT 112.120 1.720 113.170 2.570 ;
        RECT 134.470 2.010 135.070 2.570 ;
      LAYER met4 ;
        RECT 156.150 4.650 157.460 5.450 ;
        RECT 45.750 1.070 47.180 2.040 ;
        RECT 67.740 1.500 69.320 2.560 ;
        RECT 46.150 1.000 46.770 1.070 ;
        RECT 68.240 1.000 68.840 1.500 ;
        RECT 89.590 1.280 91.650 2.590 ;
        RECT 111.600 1.470 113.850 2.850 ;
        RECT 134.110 1.700 135.430 2.800 ;
        RECT 90.320 1.000 90.930 1.280 ;
        RECT 112.400 1.000 113.010 1.470 ;
        RECT 134.480 1.000 135.080 1.700 ;
        RECT 156.560 1.000 157.160 4.650 ;
        RECT 46.150 0.990 46.160 1.000 ;
        RECT 46.760 0.990 46.770 1.000 ;
        RECT 90.920 0.990 90.930 1.000 ;
  END
END tt_um_ardratag_tt_relu
END LIBRARY

